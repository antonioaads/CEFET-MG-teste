module processador_top();

wire clock;
wire []
registrador_16bits(clock, din, dout);

endmodule